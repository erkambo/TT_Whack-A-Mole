`default_nettype none

// ============================================================================
// Countdown Timer Module
// ============================================================================
module countdown_timer(
    input  wire        clk,
    input  wire        rst_n,
    input  wire        enable,
    input  wire [15:0] preset,
    output reg  [15:0] count,
    output wire        done
);
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            count <= preset;
        else if (enable && count != 16'd0)
            count <= count - 1'b1;
    end
    assign done = (count == 16'd0);
endmodule


// ============================================================================
// Round Timer Module
// ============================================================================
module round_timer(
    input  wire        clk,
    input  wire        rst_n,
    input  wire        enable,
    input  wire        reset_round,
    input  wire [15:0] preset,
    output reg  [15:0] count,
    output wire        expired
);
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n || reset_round)
            count <= preset;
        else if (enable && count != 16'd0)
            count <= count - 1'b1;
    end
    assign expired = (count == 16'd0);
endmodule


// ============================================================================
// Pattern Generator: LFSR‐based, picks exactly num_lit bits
// ============================================================================
module pattern_gen(
    input  wire        clk,
    input  wire        rst_n,
    input  wire [15:0] seed,
    input  wire [2:0]  num_lit,
    output reg  [6:0]  pattern
);
    reg [15:0] lfsr;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            lfsr <= seed;
        else
            lfsr <= {lfsr[14:0], lfsr[15]^lfsr[13]^lfsr[12]^lfsr[10]};
    end

    integer i, count;
    always @(*) begin
        pattern = 7'b0;
        count   = 0;
        for (i = 0; i < 7; i = i + 1) begin
            if (lfsr[i] && count < num_lit) begin
                pattern[i] = 1'b1;
                count = count + 1;
            end
        end
        for (i = 0; i < 7; i = i + 1) begin
            if (count < num_lit && pattern[i] == 1'b0) begin
                pattern[i] = 1'b1;
                count = count + 1;
            end
        end
    end
endmodule


// ============================================================================
// Game FSM for pattern‐pressing
// ============================================================================
module game_fsm_patterns(
    input  wire        clk,
    input  wire        rst_n,
    input  wire [6:0]  pattern,
    input  wire [7:0]  btn_sync,
    input  wire        game_end,
    input  wire        round_expired,
    output reg         reset_round,
    output reg  [7:0]  lockout,
    output reg  [7:0]  score_cnt,
    output reg  [6:0]  pattern_latched
);
    typedef enum reg { WAIT = 1'b0, NEXT = 1'b1 } state_t;
    state_t state;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            pattern_latched <= 7'b0;
            lockout         <= 8'd0;
            score_cnt       <= 8'd0;
            state           <= NEXT;
            reset_round     <= 1'b1;
        end else if (!game_end) begin
            case (state)
                NEXT: begin
                    pattern_latched <= pattern;
                    lockout         <= 8'd0;
                    reset_round     <= 1'b1;
                    state           <= WAIT;
                end

                WAIT: begin
                    reset_round <= 1'b0;
                    if ((btn_sync[6:0] & pattern_latched) == pattern_latched
                        && pattern_latched != 7'b0) begin
                        score_cnt <= score_cnt + 1;
                        state     <= NEXT;
                    end else if (|(btn_sync[6:0] & ~pattern_latched)) begin
                        lockout <= btn_sync;
                        state   <= WAIT;
                    end else if (round_expired) begin
                        state <= NEXT;
                    end
                end
            endcase
        end
    end
endmodule


// ============================================================================
// 7‐segment Driver: shows pattern or final score (lower hex digit)
// ============================================================================
module seg7_driver_patterns(
    input  wire [6:0]  pattern,
    input  wire        game_end,
    input  wire [3:0]  score_nibble,
    output reg  [6:0]  seg,
    output reg         dp
);
    always @(*) begin
        seg = ~pattern;
        dp  = 1'b1;
        if (game_end) begin
            dp = 1'b0;
            case (score_nibble)
                4'h0: seg = 7'b1000000;
                4'h1: seg = 7'b1111001;
                4'h2: seg = 7'b0100100;
                4'h3: seg = 7'b0110000;
                4'h4: seg = 7'b0011001;
                4'h5: seg = 7'b0010010;
                4'h6: seg = 7'b0000010;
                4'h7: seg = 7'b1111000;
                4'h8: seg = 7'b0000000;
                4'h9: seg = 7'b0010000;
                4'hA: seg = 7'b0001000;
                4'hB: seg = 7'b0000011;
                4'hC: seg = 7'b1000110;
                4'hD: seg = 7'b0100001;
                4'hE: seg = 7'b0000110;
                4'hF: seg = 7'b0001110;
                default: seg = 7'b1000000;
            endcase
        end
    end
endmodule


// ============================================================================
// Core game (with ena port, as requested)
// ============================================================================
module tt_um_whack_a_mole(
    input  wire        clk,
    input  wire        rst_n,
    input  wire        ena,
    input  wire [7:0]  ui_in,
    input  wire [7:0]  uio_in,
    output wire [7:0]  uo_out,
    output wire [7:0]  uio_out,
    output wire [7:0]  uio_oe,
    output wire        game_end,
    output wire        round_expired,
    output wire [7:0]  lockout
);
    wire [7:0] btn_sync        = ui_in & ~lockout;
    wire [7:0] score;
    wire [15:0] timer_count;
    wire [15:0] round_count;
    wire [6:0]  generated_pattern;
    wire        reset_round;
    wire [7:0]  fsm_lockout;

    // suppress unused uio_in warning
    wire _unused_uio = &uio_in;

    // difficulty curves
    wire [15:0] round_preset = (score <  8'd5)  ? 16'd5000 :
                               (score <  8'd10) ? 16'd4000 :
                               (score <  8'd20) ? 16'd3000 :
                                                   16'd2000;
    wire [2:0]  num_lit      = (score <  8'd5)  ? 3'd1 :
                               (score <  8'd10) ? 3'd2 :
                               (score <  8'd20) ? 3'd3 :
                                                   3'd4;

    wire [6:0] seg;
    wire       dp;

    assign lockout       = fsm_lockout;
    assign uo_out        = {dp, seg};
    assign uio_out       = score;
    assign uio_oe        = 8'hFF;

    countdown_timer timer_inst (
        .clk    (clk),
        .rst_n  (rst_n & ena),
        .enable (ena && !game_end),
        .preset (16'd60000),
        .count  (timer_count),
        .done   (game_end)
    );

    round_timer round_timer_inst (
        .clk         (clk),
        .rst_n       (rst_n & ena),
        .enable      (ena && !game_end),
        .reset_round (reset_round),
        .preset      (round_preset),
        .count       (round_count),
        .expired     (round_expired)
    );

    pattern_gen pattern_gen_inst (
        .clk     (clk),
        .rst_n   (rst_n & ena),
        .seed    (timer_count),
        .num_lit (num_lit),
        .pattern (generated_pattern)
    );

    game_fsm_patterns fsm_inst (
        .clk            (clk),
        .rst_n          (rst_n & ena),
        .pattern        (generated_pattern),
        .btn_sync       (btn_sync),
        .game_end       (game_end),
        .round_expired  (round_expired),
        .reset_round    (reset_round),
        .lockout        (fsm_lockout),
        .score_cnt      (score),
        .pattern_latched()
    );

    seg7_driver_patterns drv_inst (
        .pattern      (generated_pattern),
        .game_end     (game_end),
        .score_nibble (score[3:0]),
        .seg          (seg),
        .dp           (dp)
    );
endmodule


// ============================================================================
// Wrapper for cocotb: top‐level is 'dut', instantiates core as instance 'dut'
// ============================================================================  
module dut(
    input  wire        clk,
    input  wire        rst_n,
    input  wire [7:0]  ui_in,
    output wire [7:0]  uo_out,
    output wire [7:0]  uio_out,
    output wire [7:0]  uio_oe,
    output wire        game_end,
    output wire        round_expired,
    output wire [7:0]  lockout
);
    tt_um_whack_a_mole dut (
        .clk           (clk),
        .rst_n         (rst_n),
        .ena           (1'b1),
        .ui_in         (ui_in),
        .uio_in        (8'h00),
        .uo_out        (uo_out),
        .uio_out       (uio_out),
        .uio_oe        (uio_oe),
        .game_end      (game_end),
        .round_expired (round_expired),
        .lockout       (lockout)
    );
endmodule

`default_nettype wire
